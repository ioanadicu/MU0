// COMP12111 Exercise 3 - MU0_Alu 
// Version 2024. P W Nutter
//
// MU0 ALU design 
//
// Comments:
//
// According Table 2: ALU operations as a function of M, we implement the following cases
// M = 00 -> Y
// M = 01 -> X + Y
// M = 10 -> x + 1
// M = 11 -> X - Y (for this we'll use 2's complement to avoid substraction: invert all bits and add 1
// We will use Q for output of the function
//

// Do not touch the following line it is required for simulation 
`timescale 1ns/100ps
`default_nettype none

// module header

module MU0_Alu (
               input  wire [15:0]  X, 
               input  wire [15:0]  Y, 
               input  wire [1:0]   M, 
               output reg  [15:0]  Q
	       );

// behavioural description for the ALU

always @(*) // asynchronous (w/o global clock), combinatorial (the output depends on current inputs), we use = blocking assignment
begin
	case(M) // the operation depends on the status of the 2-bit control signal M
		2'b00:	Q = Y;	// if M is 00 output Y
		2'b01:	Q = X + Y;	// if M is 01 output X + Y
		2'b10:	Q = X + 1;	// if M is 10 output X + 1
		2'b11:	Q = X + (~Y + 1);	// if M is 11 output X - Y: we're doing the substraction using two's complement according to instructions
		default: Q = 16'bxxxx_xxxx_xxxx_xxxx; // default case for good practice
	endcase
end


endmodule 

// for simulation purposes, do not delete
`default_nettype wire
