// COMP12111 Exercise 3 - MU0_Mux12 Testbench
// Version 2024. P W Nutter
//
// Testbench for the 2-to-1 12-bit MUX
// DUT is instantiated for you.
// Need to complete the test stimulus.
//
// Comments:
//
// Testing pairs of inputs, covering unknown modes and different number combinations
// for each S input.
// 
// All unused inputs set to X.
// Xs will tend to propagate and expose faults in digital simulations
//

// Do not touch the following lines as they required for simulation 
`timescale  1ns / 100ps
`default_nettype none

module MU0_Mux12_Testbench();

//  Internal signals have been defined for you
//  and must be used for this excercise 
//  DO NOT alter the names of these signals 

reg   [11:0] A, B;
reg          S; 
wire  [11:0] Q; 


// The design has been instantiated for you below:

MU0_Mux12 top(.A(A), .B(B), .S(S), .Q(Q) );


/* Comment block

#VALUE      creates a delay of VALUE ps
a=VALUE;    sets the value of input 'a' to VALUE
$stop;      tells the simulator to stop

*/

initial
begin
// Enter you stimulus below this line
// -------------------------------------------------------

	S = 1'bx; 			// Unknown mode
	A = 12'hxxx; 	
	B = 12'hxxx; 
	// Expect Q = 12'hxxx
	
	#100;
	S = 1'b0;			// Q = A mode
	A = 12'h222;
	B = 12'hxxx;
	// Expect Q = 12'h222

	#100;
	S = 1'b1;			// Q = B mode
	A = 12'hxxx;
	B = 12'h444;
	// Expect Q = 12'h444

	#100;
	S = 1'bx; 			// Unknown mode
	A = 12'hxxx; 	
	B = 12'hxxx; 
	// Expect Q = 12'hxxx

// -------------------------------------------------------
// Please make sure your stimulus is above this line

#100 $stop;
end


endmodule

`default_nettype wire
