// COMP12111 Exercise 3 - MU0_Mux16 Testbench
// Version 2024. P W Nutter
//
// Testbench for the 2-to-1 16-bit MUX
// DUT is instantiated for you.
// Need to complete the test stimulus.
//
// Comments:
//
// Testing pairs of inputs, covering unknown modes and different number combinations
// for each S input.
// 
// All unused inputs set to X.
// Xs will tend to propagate and expose faults in digital simulations
//

// Do not touch the following lines as they required for simulation 
`timescale  1ns / 100ps
`default_nettype none

module MU0_Mux16_Testbench();

//  Internal signals have been defined for you
//  and must be used for this excercise 
//  DO NOT alter the names of these signals 

reg   [15:0] A, B;
reg          S; 
wire  [15:0] Q;


// The design has been instantiated for you below:

MU0_Mux16 top(.A(A), .B(B), .S(S), .Q(Q) );


/* Comment block

#VALUE      creates a delay of VALUE ps
a=VALUE;    sets the value of input 'a' to VALUE
$stop;      tells the simulator to stop

*/

initial
begin
// Enter you stimulus below this line
// -------------------------------------------------------

	S = 1'bx; 			// Unknown mode
	A = 16'hxxxx; 	
	B = 16'hxxxx; 
	// Expect Q = 12'hxxxx
	
	#100;
	S = 1'b0;			// Q = A mode
	A = 16'h2222;
	B = 16'hxxxx;
	// Expect Q = 12'h2222

	#100;
	S = 1'b1;			// Q = B mode
	A = 16'hxxxx;
	B = 16'h4444;
	// Expect Q = 12'h4443

	#100;
	S = 1'bx; 			// Unknown mode
	A = 16'hxxxx; 	
	B = 16'hxxxx; 
	// Expect Q = 12'hxxxx

// -------------------------------------------------------
// Please make sure your stimulus is above this line

#100 $stop;
end


endmodule

`default_nettype wire
