// COMP12111 Exercise 1 - Combinatorial Design
//
// Version 2024. P W Nutter
//
// To do:
// - produce behavioural description of the multisegment decoder
//
// DO NOT change the interface to this design 
//
// Document your code - marks may be awarded/lost for the 
// quality of the comments given. Please document in the header 
// the changes made, when and by whom.
//
// Comments:
//

`timescale  1ns / 100ps
`default_nettype none

module Display_Decoder (input wire  [3:0]  input_code,       // bcd input
			            output reg 	[14:0] segment_pattern); // segment code output

// provide Verilog that described the required behaviour of the
// combinatorial design
// -----------------------------------------------------------------







endmodule  // end of module Display_Decoder

`default_nettype wire
